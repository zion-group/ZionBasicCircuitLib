///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Use place   : ZionBasicCircuitLib_**RcDff
// Author      : Wenheng Ma
// Date        : 2019-11-05
// Version     : 1.0
// Parameter   : None
// Description :
//   This This macro definition is used in ZionBasicCircuitLib_ClrEnRcDff,
//   ZionBasicCircuitLib_ClrRcDff,ZionBasicCircuitLib_EnRcDff.
//   The macro defines the type of reset, the user can change the content of 
//   the macro definition as needed. The compilation order of this file must be 
//   before ZionBasicCircuitLib_ClrEnRcDff,ZionBasicCircuitLib_ClrRcDff,ZionBasicCircuitLib_EnRcDff. 
// Modification History:
//    Date    |   Author   |   Version   |   Change Description
//======================================================================================================================
// 2019-10-29 |  Yudi Gao  |     1.0     |   Original Version
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`define RST_CFG_SYN_HIGH 